import fidl "intf\\fidl\\com\\harman\\connectivity\\BtService.fidl"
import fidl "intf\\fidl\\com\\harman\\connectivity\\Phonebook.fidl"
import fidl "intf\\fidl\\com\\harman\\connectivity\\AndroidAutoDomainSvc.fidl"
import fidl "intf\\fidl\\com\\harman\\connectivity\\MirrorLinkDomainSvc.fidl"
import fidl "intf\\fidl\\com\\harman\\connectivity\\CarPlayDomainSvc.fidl"
import fidl "intf\\fidl\\com\\harman\\connectivity\\iAP2DevCtrl.fidl"
import fidl "intf\\fidl\\com\\harman\\connectivity\\WifiService.fidl"
import fidl "intf\\fidl\\com\\harman\\connectivity\\iAP1DevCtrl.fidl"
import cdl "../swpl/orinoco_base.cdl"
import cdl "../genivi/Genivi.cdl"
import cdl "../audio/audioManager.cdl"
import cdl "../audio/wavePlayer.cdl"


/*
 * Package delivered by CoC Connectivity for Orinoco2.0
 */
package cc_connectivity{
	generator true
	/*
	 * Bluetooth Service
	 */

	 component BTService extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.BtService as inst0
		/*
		 * PhoneBook control
		 */
		consumes interface com.harman.connectivity.PhoneBook instance dynamic as pimDbProxy
		/*
		 * Audio Management control
		 */
		provides interface org.genivi.am.routinginterface.RoutingControl as btRoutCtrl 
		consumes interface org.genivi.am.commandinterface.CommandControl instance audioManager::commandInst as commandInst
		consumes interface org.genivi.am.routinginterface.RoutingControlObserver instance audioManager::routingInst as routingInst
		/*
		 * WavePlayer control
		 */
        consumes interface com.harman.audio.waveplayer.wavePlayer instance providerComp::wavePlayerProvider as wavePlayerInst
	}
	
	component BTsvcTestClient {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.BtService instance dynamic as btProxy
		
	}
	
	/*
	 * Pim Db Service
	 */
	component PimDbService extends orinoco_component {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.PhoneBook as inst0
		/*
		 * BtService control
		 */
		consumes interface com.harman.connectivity.BtService instance dynamic as btProxy
	}
	
	component PimDbTestClient {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.PhoneBook instance dynamic as pimDbProxy
		
	}
	
	/*
	 * Carplay Service
	 */
	 component CarPlayDomainService extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.CarPlayDomainSvc as inst0
		consumes interface com.harman.connectivity.iAP2DevCtrl instance dynamic as iAP2Proxy
		/*
		* Audio Management control
		*/
		provides interface org.genivi.am.routinginterface.RoutingControl as cPlayRoutCtrl
		consumes interface org.genivi.am.commandinterface.CommandControl instance audioManager::commandInst as commandInst
		consumes interface org.genivi.am.routinginterface.RoutingControlObserver instance audioManager::routingInst as routingInst
		consumes interface com.harman.connectivity.BtService instance dynamic as btProxy
	}
	
	component cPlayTestClient {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.CarPlayDomainSvc instance dynamic as cPlayProxy
		
	}

	/*
	 * AndroidAuto Service
	 */
	component AndroidAutoDomainSvc extends orinoco_component {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.AndroidAutoDomainSvc as inst0
		/*
		 * Audio Management control
		 */
		provides interface org.genivi.am.routinginterface.RoutingControl as aAutoRoutCtrl
		consumes interface org.genivi.am.commandinterface.CommandControl instance audioManager::commandInst as commandInst
		consumes interface org.genivi.am.routinginterface.RoutingControlObserver instance audioManager::routingInst as routingInst
		consumes interface com.harman.connectivity.BtService instance dynamic as btProxy
	}
	
	component androidAutoTestClient {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.AndroidAutoDomainSvc instance dynamic as androidAutoProxy
		
	}

	/*
	* MirrorLink Service
	*/	
	component MirrorLinkDomainSvc extends orinoco_component {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.MirrorLinkDomainSvc as inst0
		/*
		 * Audio Management control
		 */
		provides interface org.genivi.am.routinginterface.RoutingControl as mLinkRoutCtrl
		consumes interface org.genivi.am.commandinterface.CommandControl instance audioManager::commandInst as commandInst
		consumes interface org.genivi.am.routinginterface.RoutingControlObserver instance audioManager::routingInst as routingInst
	}
	
	component mLinkTestClient {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.MirrorLinkDomainSvc instance dynamic as mLinkProxy
		
	}
	
	/*
	* IAP2 Service
	*/	
	component iAP2DevCtrl extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.iAP2DevCtrl as inst0
		
	}
	component iAP2DevCtrlTest {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.iAP2DevCtrl instance dynamic as iAP2Proxy
	}
    
    /*
	* IAP1 Service
	*/	
	component iAP1DevCtrl extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.iAP1DevCtrl as inst0
		
	}
	component iAP1DevCtrlTest {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.iAP1DevCtrl instance dynamic as iAP1Proxy
	}
    
	/*
	 * Wi-Fi Service
	 */
	component WifiService extends orinoco_component {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.connectivity.WifiService as inst0
	}
	
	component WifiServiceTestClient {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.connectivity.WifiService instance dynamic as wlanProxy
		
	}	

}