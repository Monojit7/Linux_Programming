import fidl "intf\\fidl\\com\\harman\\RVCservice\\RVCClient.fidl"

/*
 * Package delivered by CoC Platform Software for Orinoco2.0
 */
package RVCClient{
	generator true

	component RVCService	{
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.RVCservice.RVC as inst0
	}
	
	component RVCServiceTest	{
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.RVCservice.RVC instance RVCService::inst0 as RVCProxy
	}
}

