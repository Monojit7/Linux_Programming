import fidl "./intf/fidl/com/harman/audio/ecnr.fidl"

import cdl "../swpl/orinoco_base.cdl"

/*
 * 
 */ 


package cc_audio{
	generator true
	
	component ecnr extends orinoco_component {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.audio.ecnr.ecnr as ecnrInst
	}
	
	component ecnrClient {
		buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.audio.ecnr.ecnr instance ecnr::ecnrInst as ecnrProxy
	}
}