
import cdl "cc_swpl.cdl"
import cdl "../../packages/connectivity/cc_connectivity.cdl"

import fidl "intf/fidl/com/harman/swdl/SoftwareDownload.fidl"

package orinoco_platform_swdl {
	generator true
		
		component SoftwareDownload{
			buildType CMake
			language cpp
			rpc dbus
			provides interface com.harman.swdl.SoftwareDownload as swdl 
			consumes interface org.genivi.NodeStateManager.Consumer instance NodeStateManager::inst0 as nsm_consumer 	
			consumes interface org.genivi.NodeStateManager.LifecycleControl instance NodeStateManager::inst1 as proxyInst		
			consumes interface com.harman.connectivity.WifiService instance dynamic as wlanProxy
			consumes interface com.harman.connectivity.WifiService instance WifiService::inst0 as wlanProxy
		}
}
