import fidl "intf/fidl/com/harman/tuner/OrinocoTuner.fidl"
import fidl "../genivi/intf/fidl/org/genivi/am/RoutingInterface.fidl"
import cdl "../swpl/orinoco_base.cdl"
import cdl "../audio/audioManager.cdl"

/*
 * Package delivered by CoC Tuner for Orinoco2.0
 */
package cc_tuner{
	
	generator true

	component TunerApp extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.tuner.OrinocoTuner as inst0
		provides interface org.genivi.am.routinginterface.RoutingControl as inst0
		consumes interface org.genivi.am.routinginterface.RoutingControlObserver instance audioManager::routingInst as routingInst
	}
	
	component TunerAppTest {
	 	buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.tuner.OrinocoTuner instance TunerApp::inst0 as OrinocoTunerProxy
	}
}