//Import the base orinoco component
import cdl "packages/swpl/orinoco_base.cdl"
import cdl "packages/media/cc_media.cdl"

package oakland_mmpres{
	generator true
	
	component mpres extends orinoco_component{
		buildType CMake
		language cpp
		rpc dbus
		
		
		/*
		 * MediaOne
		 */
		consumes interface org.genivi.mediamanager.Browser instance MediaOneService::inst0 as mediaBrowser
		consumes interface org.genivi.mediamanager.Indexer instance MediaOneService::inst0 as mediaIndexer
		consumes interface org.genivi.mediamanager.Player instance MediaOneService::inst0 as mediaPlayer
		consumes interface com.harman.media.DeviceManager instance MediaOneService::inst0 as deviceManager
		consumes interface com.harman.media.PlayerExt instance MediaOneService::inst0 as playerExt
		consumes interface com.harman.media.ImageProcess instance ImageService::inst0 as imageProc
		
				
	}
}