import fidl "../genivi/intf/fidl/org/genivi/NodeStateManager/Consumer.fidl"
import cdl "cc_swpl.cdl"

package orinoco_base{

generator true
	/*
	 * 	Every Orinoco component shall derive from the orinoco component.
 	 */	
    contains package cc_swpl
	abstract component orinoco_component
	{
		consumes interface org.genivi.NodeStateManager.Consumer instance NodeStateManager::inst0 as nsm_consumer 
	}

}




