import fidl "intf\\fidl\\com\\harman\\media\\BaseType.fidl"
import fidl "intf\\fidl\\com\\harman\\media\\DeviceManager.fidl"
import fidl "intf\\fidl\\com\\harman\\media\\PlayerExt.fidl"
import fidl "intf\\fidl\\com\\harman\\media\\ImageProcess.fidl"
import fidl "intf\\fidl\\com\\harman\\media\\MediaSetting.fidl"

import cdl "../swpl/orinoco_base.cdl"
import cdl "../genivi/Genivi.cdl"
import cdl "../connectivity/cc_connectivity.cdl"
import cdl "../audio/audioManager.cdl"

using package orinoco_base

/*
 * Package delivered by CoC Media for Orinoco2.0
 */
package cc_media{
	generator true
	
	/*
	 * MediaOne Service
	 */
	 component MediaOneService extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.media.DeviceManager as inst0
		provides interface com.harman.media.PlayerExt as inst0
		provides interface com.harman.media.MediaSetting as inst0
		provides interface org.genivi.mediamanager.Browser as inst0
		provides interface org.genivi.mediamanager.Indexer as inst0
		provides interface org.genivi.mediamanager.Player as inst0
		provides interface org.genivi.am.routinginterface.RoutingControl as Inst
		
		consumes interface com.harman.connectivity.iAP2DevCtrl instance dynamic as iAP2Proxy
		consumes interface org.genivi.am.routinginterface.RoutingControlObserver instance audioManager::routingInst as RoutingControlObserverProxy
	}
	
	component mediaone_client extends orinoco_component {
		buildType CMake
		language cpp
		rpc dbus
		
		consumes interface com.harman.media.DeviceManager instance MediaOneService::inst0 as dmProxy
		consumes interface com.harman.media.PlayerExt instance MediaOneService::inst0 as peProxy
		consumes interface org.genivi.mediamanager.Browser instance MediaOneService::inst0 as brProxy
		consumes interface org.genivi.mediamanager.Indexer instance MediaOneService::inst0 as idProxy
		consumes interface org.genivi.mediamanager.Player instance MediaOneService::inst0 as plProxy
	}
	
	component ImageService extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.media.ImageProcess as inst0
	}
	
	component ImageService_client extends orinoco_component {
	 	buildType CMake
		language cpp
		rpc dbus
		consumes interface com.harman.media.ImageProcess instance ImageService::inst0 as isProxy
	}
	
}