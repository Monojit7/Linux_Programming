//Import the base orinoco component
import cdl "packages/swpl/orinoco_base.cdl"

//Import cdls
import cdl 'packages/connectivity/cc_connectivity.cdl'
import cdl "packages/genivi/Genivi.cdl"
import cdl "packages/tuner/cc_tuner.cdl"
import cdl "packages/audio/audioManager.cdl"
import cdl "packages/connectivity/CarLifeDomainSvc.cdl"
import cdl "packages/media/cc_media.cdl"
//import cdl "packages/swpl/orinoco_swdl.cdl"
import fidl "packages/swdl/SoftwareDownload.fidl"

//Navigation fidls.. not in package format !
import fidl "packages/nav/ctrl/mapv/MapViewControl.fidl"
import fidl "packages/nav/ctrl/common/CommonTypes.fidl"
import fidl "packages/nav/ctrl/configuration/Configuration.fidl"
import fidl "packages/nav/ctrl/configuration/ConfigurationBase.fidl"
import fidl "packages/nav/ctrl/di/LocationInput.fidl"
import fidl "packages/nav/ctrl/di/OneBoxSearch.fidl"
import fidl "packages/nav/ctrl/di/POISearch.fidl"
import fidl "packages/nav/ctrl/di/SpeechLocationInput.fidl"
import fidl "packages/nav/ctrl/di/SpeechPoiSearch.fidl"
import fidl "packages/nav/ctrl/pos/Positioning.fidl"
import fidl "packages/nav/ctrl/sim/Simulation.fidl"
import fidl "packages/nav/ctrl/icon/IconProvider.fidl"
import fidl "packages/nav/ctrl/icon/IconProvider.fidl"
import fidl "packages/nav/ctrl/common/list/ListViewBase.fidl"



package oakland_hmi{
	generator true
	
	component hmi extends orinoco_component{
		buildType CMake
		language cpp
		rpc dbus
	
		/*
		 * Telephony
		 */
		 consumes interface com.harman.connectivity.PhoneBook instance dynamic as inst0
		 consumes interface com.harman.connectivity.BtService instance dynamic as bt

		/*
		 * Projection modes
		 */
		consumes interface com.harman.connectivity.CarPlayDomainSvc instance CarPlayDomainService::inst0 as cPlayProxy
		consumes interface com.harman.connectivity.AndroidAutoDomainSvc instance AndroidAutoDomainSvc::inst0 as aAutoProxy
		consumes interface com.harman.connectivity.MirrorLinkDomainSvc instance MirrorLinkDomainSvc::inst0 as mLinkProxy
		consumes interface com.harman.service.CarLifeDomainSvc instance CarLife::inst0 as carLifeProxy

		/*
		 * Wifi  
		 */
		 consumes interface com.harman.connectivity.WifiService instance WifiService::inst0 as wlanProxy
		 				
		/*
		 * Radio
		 */
		consumes interface IVIRadio.Station.Station instance dynamic as inst0
        consumes interface IVIRadio.Configuration.Configuration instance dynamic as tunerConfig
		consumes interface IVIRadio.AdditionalService.AdditionalService instance dynamic as radioAdditionalConfig
		
		consumes interface com.harman.tuner.OrinocoTuner instance dynamic as inst0
		
		
		
		/*
		 * Audio Management control
		 */
		consumes interface org.genivi.am.commandinterface.CommandControl instance audioManager::commandInst as commandInst
		consumes interface org.genivi.am.routinginterface.RoutingControlObserver instance audioManager::routingInst as 	routingInst

		/*
		 * MediaOne
		 */
		consumes interface org.genivi.mediamanager.Browser instance MediaOneService::inst0 as mediaBrowser
		consumes interface org.genivi.mediamanager.Indexer instance MediaOneService::inst0 as mediaIndexer
		consumes interface org.genivi.mediamanager.Player instance MediaOneService::inst0 as mediaPlayer
		consumes interface com.harman.media.DeviceManager instance MediaOneService::inst0 as deviceManager
		consumes interface com.harman.media.PlayerExt instance MediaOneService::inst0 as playerExt
		consumes interface com.harman.media.ImageProcess instance ImageService::inst0 as imageProc
		
		/* 
		 * Software download for qt hmi 
		 */	
		consumes interface com.harman.swdl.SoftwareDownload instance dynamic as swdl
		
		
		
		/* Navigation***********************************************************************
         */
          /**
         * MapView
         */
        consumes interface org.harman.nav.ctrl.mapv.MapViewControl instance dynamic as MapViewControl
        
         /**
         * Configuration
         */
        consumes interface org.harman.nav.ctrl.configuration.Configuration instance dynamic as Configuration	  
        consumes interface org.harman.nav.ctrl.configuration.ConfigurationBase instance dynamic as ConfigurationBase
        
         /**
         * Location Search
         */
        consumes interface org.harman.nav.ctrl.di.LocationInput instance dynamic as LocationInput	  
        consumes interface org.harman.nav.ctrl.di.OneBoxSearch instance dynamic as OneBoxSearch
        consumes interface org.harman.nav.ctrl.di.LocationInput instance dynamic as POISearch
        consumes interface org.harman.nav.ctrl.di.LocationInput instance dynamic as SpeechLocationInput
        consumes interface org.harman.nav.ctrl.di.LocationInput instance dynamic as SpeechPoiSearch
         /**
         * icon
         */
        consumes interface org.harman.nav.ctrl.icon.IconProvider instance dynamic as IconProvider	  
        
         /**
         * Positioning
         */
        consumes interface org.harman.nav.ctrl.Positioning instance dynamic as Positioning	  
        
         /**
         * Simulation
         */
        consumes interface org.harman.nav.ctrl.Simulation instance dynamic as Simulation	  
        
        /**
         * List
         */
        consumes interface org.harman.nav.ctrl.common.list.ListViewBase instance dynamic as ListViewBase
		
	}
}