import fidl "fidl/BluetoothTypes.fidl"
import fidl "fidl/ConnectionManager.fidl"
import fidl "fidl/CallManager.fidl"
import fidl "fidl/PimDbHandler.fidl"

import cdl "../connectivity/cc_connectivity.cdl"

package btpres{
	generator true

	component btpres
	{
		buildType CMake
		language cpp
		rpc dbus

		provides interface com.harman.btpres.ConnectionManager as connectionManager
		provides interface com.harman.btpres.CallManager as callManager
		provides interface com.harman.btpres.PimDbHandler as pimManager
		
		/*
		 * BtService and PimService
		 */
		consumes interface com.harman.connectivity.BtService instance dynamic as BtServiceProxy
		consumes interface com.harman.connectivity.PhoneBook instance dynamic as PimDbProxy
	}

	component btprestest
	{
		buildType CMake
		language cpp
		rpc dbus
		
		consumes interface com.harman.btpres.ConnectionManager instance btpres::connectionManager as btpres
		consumes interface com.harman.btpres.CallManager instance btpres::callManager as btpres
		consumes interface com.harman.btpres.PimDbHandler instance btpres::pimManager as btpres
	}
}