import fidl "intf/fidl/com/harman/audio/waveplayer/wavePlayer.fidl"

package wavePlayer{
    generator true
    component providerComp  {
        language cpp
        buildType CMake
        rpc dbus
        provides interface com.harman.audio.waveplayer.wavePlayer as wavePlayerProvider
    }
     
    component consumerComp{
        language cpp
        buildType CMake
        rpc dbus
        consumes interface com.harman.audio.waveplayer.wavePlayer instance providerComp::wavePlayerProvider as wavePlayerConsumer
    }
}