import fidl "../genivi/intf/fidl/org/genivi/NodeStateManager/Consumer.fidl"
import fidl "../genivi/intf/fidl/org/genivi/NodeStateManager/LifeCycleControl.fidl"
import fidl "../genivi/intf/fidl/org/genivi/NodeStartupController1/NodeStartupController.fidl"
import fidl "../genivi/intf/fidl/org/genivi/NodeHealthMonitor/Info.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/BodyControlStatusProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/ButtonStatusProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/KeyStatusProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/PowerModeStatusProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/PulseCounterUpdateProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/TimeDateProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/VehicleSpeedProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/VINProvider.fidl"
import fidl "intf/fidl/com/harman/vehiclebroker/OperationalModeStatusProvider.fidl" 
import fidl "intf/fidl/com/harman/vehiclebroker/OrinocoSpecificData.fidl" 
import fidl "intf/fidl/com/harman/vehiclebroker/HudData.fidl" 
import fidl "intf/fidl/com/harman/pathology/Pathology.fidl"

import fidl "intf/fidl/com/harman/infotainment/systeminfrastructure/versionmanager/VersionManager.fidl"
/*
 * Packages delivered by CC_Software platform
 */
package cc_swpl{
    generator true

	/*
	 * NodeStateManager : 
	 * The node state management is the central function for information regarding the current running state of the embedded system. 
	 * The node state management also provides shutdown management, so one part of the information which is provided is the shutdown request notification to the consumers.
	 * The node state management is the last/highest level of escalation on the node and will therefore command the reset and supply control logic.
	 */
	 
	component NodeStateManager {
		buildType CMake
		language cpp
		rpc dbus
		provides interface org.genivi.NodeStateManager.Consumer as inst0
		provides interface org.genivi.NodeStateManager.LifecycleControl as inst1
	}
	
	/*
	 * Last User Context (LUC) Management
	 * Target Startup Monitoring
	 */
	component NodeStartupController {
		buildType CMake
		language cpp
		rpc dbus
		provides interface org.genivi.NodeStartupController1.NodeStartupController as inst0
	}
	/*
	 * The Node Health Monitor will work in conjunction with systemd to monitor component failures in the system.
	 * It will be responsible for :
	 * monitoring systemd to automatically record and track failures per component (i.e. application, service)
	 * providing an interface with which components can register failures when not using the systemd monitoring
	 * maintaining failure statistics over multiple lifecycles for the system and components (the service name will be used to identify and track component failures)
	 * maintaining statistics on number of failures in number of lifecycles (i.e. 3 failures in last 32 lifecycles)
	 * monitoring the wakeup and shutdown events to catch unexpected system restarts
	 */
	component NodeHealthMonitor {
		buildType CMake
		language cpp
		rpc dbus
		provides interface org.genivi.NodeHealthMonitor.Info as inst0
	}

	/*
	 * Provides interface to publish the vehicle network data (e.g. CAN)
	 */
	component VehicleDataProvider {

		language cpp
		buildType CMake
		rpc dbus
		
		provides interface com.harman.vehicle.BodyControlStatusProvider as BodyControlStatusProvider
		provides interface com.harman.vehicle.ButtonStatusProvider as ButtonStatusProvider
		provides interface com.harman.vehicle.KeyStatusProvider as KeyStatusProvider
		provides interface com.harman.vehicle.PowerModeStatusProvider as PowerModeStatusProvider
		provides interface com.harman.vehicle.PulseCounterUpdateProvider as PulseCounterUpdateProvider
		provides interface com.harman.vehicle.TimeDateProvider as TimeDateProvider
		provides interface com.harman.vehicle.VehicleSpeedProvider as VehicleSpeedProvider
		provides interface com.harman.vehicle.VINProvider as VINProvider
		provides interface com.harman.vehicle.OperationalModeStatusProvider as OperationalModeStatusProvider 
		provides interface com.harman.vehicle.HudData as HudData
		provides interface com.harman.vehicle.OrinocoSpecificData as OrinocoSpecificData
	}
 
 	/*
	* pathology is system resource monitoring component that will run for entire life cycle of the system
	* It will monitor system CPU and RAM, process CPU and RAM, process core-dump, etc
	* Also pathology will listen to systemd watchdog warning. The commonAPI interfaces will
	* be used to get the data out of pathology and provide certain tiggers as input to patholgy.
	*/
	component pathologyProvider	{
		language cpp
		buildType  CMake
		rpc dbus
		provides interface com.harman.pathology.SystemInformation as int0  
		provides interface  com.harman.pathology.TriggersToPathology as int1
	}
	
    /*
	 * Last User Context (LUC) Management
	 * Target Startup Monitoring
	 */
	component VersionManager {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.infotainment.systeminfrastructure.versionmanager.versionmanager.VersionManager as inst0
	}
 
 	/*
	 * Interface Internal to persistency and SWDL 
	 * e.g. to setup persistency data during SWDL  
	 * 
	 * -UNDER WORK-
	 */
 /*
	component PersistencyAdminService {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.persistence.Administration as inst0
	}
 */
 
 	/*
	 * -UNDER WORK-
	 */
 /*
	component RVC {
		buildType CMake
		language cpp
		rpc dbus
		provides interface com.harman.RearViewCamera as inst0
	}
 */
}

